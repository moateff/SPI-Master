`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/18/2024 03:44:18 PM
// Design Name: 
// Module Name: SPI_Master
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
//
// Description: SPI (Serial Peripheral Interface) Master
//              Creates master based on input configuration.
//              Sends a byte one bit at a time on MOSI
//              Will also receive byte data one bit at a time on MISO.
//              Any data on input byte will be shipped out on MOSI.
//
//              To kick-off transaction, user must pulse tx_start.
//              This module supports multi-byte transmissions by pulsing
//              tx_start and loading up din when ready is high.
//
//              This module is only responsible for controlling Clk, MOSI, 
//              and MISO.  If the SPI peripheral requires a chip-select, 
//              this must be done at a higher level.
//
// SPI_MODE, can be 0, 1, 2, or 3.  See above.
// Can be configured in one of 4 modes:
//              Mode | Clock Polarity (CPOL/CKP) | Clock Phase (CPHA)
//               0   |             0             |        0
//               1   |             0             |        1
//               2   |             1             |        0
//               3   |             1             |        1

module SPI_Master 
#(  
    parameter FRAME_WIDTH    = 8,         // Width of the data to be transmitted/received
              CLKS_PER_HALF  = 2          // Clock divider to control the SPI clock frequency
)(
    input  logic                     clk,        // System clock input
    input  logic                     reset,      // Reset signal to reset the SPI Master state
    input  logic [1:0]               mode,       // SPI mode: 0, 1, 2, or 3 for clock polarity (CPOL) and phase (CPHA)
    
    // TX (MOSI) Signals
    input  logic [FRAME_WIDTH - 1:0] din,        // Data to be transmitted (sent from Master to Slave)
    input  logic                     tx_start,   // Transmission start signal, triggers the data transfer
    output logic                     tx_ready,   // Indicates that SPI is ready to transmit new data
    
    // RX (MISO) Signals
    output logic [FRAME_WIDTH - 1:0] dout,       // Data received from the slave (Master In Slave Out)
    output logic                     rx_done,    // Indicates that the reception of data is done
    
    // SPI Interface
    input  logic                     miso,       // Slave-to-master data line (MISO: Master In Slave Out)
    output logic                     mosi,       // Master-to-slave data line (MOSI: Master Out Slave In)
    output logic                     sclk        // SPI clock, generated by the Master
    );

    logic cpol, cpha;

    // CPHA: Clock Phase
    // CPHA=0 means the "out" side changes the data on trailing edge of clock
    // the "in" side captures data on leading edge of clock
    // CPHA=1 means the "out" side changes the data on leading edge of clock
    // the "in" side captures data on the trailing edge of clock
    assign cpha     = mode[0];

    // CPOL: Clock Polarity
    // CPOL=0 means clock idles at 0, leading edge is rising edge.
    // CPOL=1 means clock idles at 1, leading edge is falling edge.
    assign cpol     = mode[1];
    
    typedef enum {IDLE, CPHA_DELAY, P0, P1} state_type;
    state_type state_next, state_reg;
    
    // Counter to generate the SPI clock. 
    // c_reg counts clock cycles and is used to divide the system clock 
    // to create the correct SPI clock (sclk) frequency.
    logic [$clog2(CLKS_PER_HALF * 2) - 1:0] c_next, c_reg;
    
    // Tracks the number of bits sent/received during a transaction. 
    // It ensures the correct number of bits (defined by DATA_WIDTH) are transmitted.
    logic [$clog2(FRAME_WIDTH) - 1:0]       n_next, n_reg;
    
    // Register to hold the data being transmitted. 
    // tx_reg holds the current data word and shifts bits out on the MOSI line.
    logic [FRAME_WIDTH - 1:0]               tx_next, tx_reg;
    
    // Register to store the data received from the slave on the MISO line. 
    // Data is shifted in as it arrives, and rx_reg holds the full data word once the transfer is complete.
    logic [FRAME_WIDTH - 1:0]               rx_next, rx_reg;
    
    // These registers handle the generation of the SPI clock signal (sclk). 
    // sclk_reg holds the current state of the clock, and sclk_next determines the next clock state.
    logic                                   sclk_next, sclk_reg;
    
    // w_clk is an intermediate signal used to calculate the SPI clock based on the CPHA value.
    // It helps determine when to toggle the SPI clock (sclk).
    logic                                   w_clk;

    always_ff @(posedge clk or posedge reset)
    begin
        if(reset)
        begin
            // On reset, the SPI master returns to the IDLE state, 
            // and all counters, data registers, and the SPI clock are reset.
            state_reg <= IDLE;
            c_reg     <= 0;
            n_reg     <= 0;
            tx_reg    <= 0;
            rx_reg    <= 0;
            sclk_reg  <= cpol; // Set the clock polarity based on the CPOL parameter.
        end
        else
        begin
            // On each clock cycle, update the current state and registers
            // with the next state and next register values.
            state_reg <= state_next;
            c_reg     <= c_next;
            n_reg     <= n_next;
            tx_reg    <= tx_next;
            rx_reg    <= rx_next;
            sclk_reg  <= sclk_next;
        end
    end
    
    always_comb
    begin
        // By default, set the next state to the current state, and keep the 
        // existing values for all other signals unless explicitly changed below.
        state_next    = state_reg;
        tx_ready      = 0;          // Indicates whether the SPI Master is ready to transmit data.
        rx_done       = 0;          // Signals when the data reception is complete.
        tx_next       = tx_reg;     // Default next value of tx_reg is the current tx_reg (data to be transmitted).
        rx_next       = rx_reg;     // Default next value of rx_reg is the current rx_reg (received data).
        n_next        = n_reg;      // Default next bit counter is the current value.
        c_next        = c_reg;      // Default next clock counter is the current value.

        case(state_reg)
            IDLE:
            begin
                tx_ready = 1;  // SPI Master is ready to load new data for transmission.
                
                // If a transmission start signal is detected, prepare for transmission.
                if(tx_start)
                begin
                    n_next = 0;        // Reset the bit counter for a new transmission.
                    c_next = 0;        // Reset the clock cycle counter.
                    tx_next = din;     // Load the input data (din) into the tx register for transmission.
                    state_next = P0;   // Move to the first phase (P0) of the SPI communication.
                end
            end

            P0:
            begin
                // When the clock counter reaches half the SPI clock cycle (CLKS_PER_HALF),
                // it's time to sample incoming data on the MISO line and prepare the next transmission bit.
                if(c_reg == CLKS_PER_HALF - 1)
                begin
                    c_next = 0;                   // Reset the clock cycle counter for the next phase.
                    rx_next = rx_reg << 1;        // Shift the current received bits to make room for the next incoming bit.
                    rx_next[0] = miso;            // Sample the incoming bit from the MISO line.
                    state_next = P1;              // Move to the second phase (P1) of SPI communication.
                end
                else
                    c_next = c_reg + 1;           // Otherwise, increment the clock cycle counter.
            end

            P1:
            begin
                // Similar to the P0 state, we wait until the clock counter reaches CLKS_PER_HALF.
                if(c_reg == CLKS_PER_HALF - 1)
                begin
                    // If all bits have been transmitted and received (n_reg equals DATA_WIDTH - 1),
                    // signal that the data reception is complete and go back to the IDLE state.
                    if(n_reg == FRAME_WIDTH - 1)
                    begin
                        rx_done = 1;               // Reception is complete, signal this with rx_done.
                        state_next = IDLE;         // Transition back to the IDLE state.
                    end
                    else
                    begin
                        // Otherwise, continue shifting data.
                        c_next = 0;                // Reset the clock cycle counter.
                        n_next = n_reg + 1;        // Increment the bit counter to transmit the next bit.
                        tx_next = tx_reg << 1;     // Shift the transmit data to the next bit.
                        tx_next[0] = 1'b0;         // Optionally, send a 0 as the LSB.
                        state_next = P0;           // Go back to P0 for the next bit.
                    end
                end
                else
                    c_next = c_reg + 1;            // Increment the clock cycle counter.
            end
        endcase

    end
    
    // Generate the SPI clock (sclk) based on the state and CPHA (clock phase).
    // In SPI mode 0, sclk should toggle between P0 and P1.
    // The polarity of the clock is determined by CPOL.
    assign w_clk = ((state_next == P1) && ~cpha) || ((state_next == P0) && cpha);
    
    // Depending on the clock polarity (CPOL), invert the clock signal if CPOL is 1.
    assign sclk_next = cpol ? ~w_clk : w_clk;
    
    // Assign the registered clock signal (sclk_reg) to the output sclk.
    assign sclk = sclk_reg;

    // The MOSI line outputs the most significant bit of the transmit register (tx_reg).
    // If the state is IDLE, MOSI is not transmitting, so it defaults to 'x' (unknown).
    assign mosi = (state_reg == IDLE) ? 1'bx : tx_reg [FRAME_WIDTH - 1];
    
    // Assign dout (output data) to rx_reg when rx_done is high, indicating a full word has been received.
    assign dout = rx_done ? rx_reg : dout;

    
endmodule
